library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Package Declaration Section
package theta_control_pkg is

    type phase_arr is array (integer range<>) of std_logic_vector(31 downto 0);
 
   
end package theta_control_pkg;
 
-- Package Body Section
--package body theta_control_pkg is
 
 
--end package body theta_control_pkg;
